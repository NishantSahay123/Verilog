module anddelay(input a,b, output c);
and #(4) and_gate_2(c,a,b);
endmodule