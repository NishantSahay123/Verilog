module and_or_xor_gate(input a,b, output c,d,e);
and(c, a, b);
or(d, a, b);
xor(e, a, b);
endmodule